library verilog;
use verilog.vl_types.all;
entity inputdev is
    port(
        din             : in     vl_logic_vector(31 downto 0);
        dout            : out    vl_logic_vector(31 downto 0)
    );
end inputdev;
